`timescale 1ns / 1ps

module my_FPHUB_adder #(
    parameter int M = 23,              // Mantissa size
    parameter int E = 8,               // Exponent size
    parameter int special_case = 7,    // Number of special cases (including non-special)
    // Parameters for mantissa extension:
    parameter int sign_mantissa_bit  = 1,
    parameter int one_implicit_bit   = 1,
    parameter int ilsb_bit           = 1,
    parameter int extra_bits_mantissa = 1 + sign_mantissa_bit + one_implicit_bit + ilsb_bit
)(
    input  logic start,             // Start signal
    input  logic signed [E+M:0] X,  // Input X
    input  logic signed [E+M:0] Y,  // Input Y
    output logic finish,            // Finish signal
    output logic [E+M:0] Z          // Output Z
);

// Test numbers
logic [E+M:0] X_prueba, Y_prueba;
assign X_prueba = 9'b011110011;
assign Y_prueba = 9'b111111000;

//--------------------------------------------------------------------------------------------------
// Special case identification
//--------------------------------------------------------------------------------------------------
logic [M+E:0] special_result;
logic [$clog2(special_case)-1:0] X_special_case, Y_special_case;
logic special_case_detected;

special_cases_detector #(E, M, special_case) special_cases_inst (
    .X(X),
    .Y(Y),
    .X_special_case(X_special_case),
    .Y_special_case(Y_special_case)
);

special_result_for_adder #(E, M, special_case) special_result_inst (
    .X(X),
    .Y(Y),
    .X_special_case(X_special_case),
    .Y_special_case(Y_special_case),
    .special_result(special_result)
);

//--------------------------------------------------------------------------------------------------
// Exponent difference calculation
//--------------------------------------------------------------------------------------------------
logic signed [E:0] diff;
logic [E:0] diff_abs;
logic X_greater_than_Y;
logic Ex_equal_Ey;

Exponent_difference #(E) Exponent_difference_inst (
    .Ex(X[E+M-1:M]),
    .Ey(Y[E+M-1:M]),
    .dif(diff),
    .X_greater_than_Y(X_greater_than_Y),
    .Ex_equal_Ey(Ex_equal_Ey)
);

//--------------------------------------------------------------------------------------------------
// Determination of effective operation and result sign
//--------------------------------------------------------------------------------------------------
logic subtraction, Sz;
assign subtraction = X[E+M] ^ Y[E+M];

//--------------------------------------------------------------------------------------------------
// Mantissa and sign organization
//--------------------------------------------------------------------------------------------------
// Internal signals defined with width M+extra_bits_mantissa
logic signed [M+extra_bits_mantissa-1:0] M_major, M_minor, M_minor_ready;
logic [E-1:0] Ez;
// Flag indicating other modules should print values
logic print;
// ILSB bits
logic ilsb_x, ilsb_y;

//--------------------------------------------------------------------------------------------------
// Alignment of the smaller mantissa using a wire
//--------------------------------------------------------------------------------------------------
logic [M+extra_bits_mantissa-1:0] M_minor_aligned;

shifter #(
  .M(M),
  .E(E),
  .extra_bits_mantissa(extra_bits_mantissa)
) shifter_inst (
  .number_input(M_minor_ready),
  .shift_amount(diff_abs),
  .right_shift(1'b1),
  .arithmetic_shift(1'b1),
  .number_output(M_minor_aligned),
  .print(print)
);

//--------------------------------------------------------------------------------------------------
// Mantissa Addition/Subtraction
//--------------------------------------------------------------------------------------------------
logic signed [M+extra_bits_mantissa-1:0] M_result, M_result_ready, M_normalize;

logic [$clog2(M+extra_bits_mantissa-sign_mantissa_bit-1):0] shift_LZA;
logic [E:0] Ez_normalized;
logic [E+M:0] result;

LZD #(
      .M(M),
      .extra_bits_mantissa(extra_bits_mantissa),
      .sign_mantissa_bit(sign_mantissa_bit)
) LZA_inst (
      .A(M_result_ready[M+extra_bits_mantissa-sign_mantissa_bit-1:0]),
      .shift_amt(shift_LZA),
      .print(print)
);
always_comb begin
    if (start) begin
        // Determine the sign of the result
        Sz = (X_greater_than_Y) ? X[E+M] : Y[E+M];

        // Define ILSB for special cases (default always 1)
        ilsb_x = (X_special_case == 5 || X_special_case == 6) ? 1'b0 : 1'b1;
        ilsb_y = (Y_special_case == 5 || Y_special_case == 6) ? 1'b0 : 1'b1;

        // Assign major and minor mantissas
        M_major = (X_greater_than_Y) ? 
            { {sign_mantissa_bit{1'b0}}, {one_implicit_bit{1'b1}}, X[M-1:0], ilsb_x,
            {(extra_bits_mantissa - (sign_mantissa_bit+one_implicit_bit+ilsb_bit)){1'b0} } } :
            { {sign_mantissa_bit{1'b0}}, {one_implicit_bit{1'b1}}, Y[M-1:0], ilsb_y,
            {(extra_bits_mantissa - (sign_mantissa_bit+one_implicit_bit+ilsb_bit)){1'b0} } };

        M_minor = (X_greater_than_Y) ? 
            { {sign_mantissa_bit{1'b0}}, {one_implicit_bit{1'b1}}, Y[M-1:0], ilsb_y,
            {(extra_bits_mantissa - (sign_mantissa_bit+one_implicit_bit+ilsb_bit)){1'b0} } } :
            { {sign_mantissa_bit{1'b0}}, {one_implicit_bit{1'b1}}, X[M-1:0], ilsb_x,
            {(extra_bits_mantissa - (sign_mantissa_bit+one_implicit_bit+ilsb_bit)){1'b0} } };

        // The output exponent is the largest of the two unless normalization is needed
        Ez = (X_greater_than_Y) ? X[E+M-1:M] : Y[E+M-1:M];

        // Flag for special cases (specifically zero and infinity cases)
        if ((X_special_case >= 1 && X_special_case <= 4) || (Y_special_case >= 1 && Y_special_case <= 4))
            special_case_detected = 1;
        else
            special_case_detected = 0;

        // Calculate absolute value of exponent difference
        diff_abs = (diff < 0) ? -diff : diff;

        // Remaining comments are translated similarly (truncated here due to length limitations)

    end
end

assign Z = (special_case_detected) ? special_result : result;
assign finish = 1'b1; // Indicate that operation has finished

endmodule